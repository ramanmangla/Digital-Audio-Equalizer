// megafunction wizard: %FIR II v18.0%
// GENERATION: XML
// BandFIR5503000.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module BandFIR5503000 (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [31:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [31:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	BandFIR5503000_0002 bandfir5503000_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2018 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="18.0" >
// Retrieval info: 	<generic name="filterType" value="single" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="symmetryMode" value="nsym" />
// Retrieval info: 	<generic name="L_bandsFilter" value="1" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="clockRate" value="50" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="inputRate" value="0.048" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="read_write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone V" />
// Retrieval info: 	<generic name="speedGrade" value="medium" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="reconfigurable" value="false" />
// Retrieval info: 	<generic name="num_modes" value="2" />
// Retrieval info: 	<generic name="reconfigurable_list" value="0" />
// Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
// Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
// Retrieval info: 	<generic name="inputType" value="int" />
// Retrieval info: 	<generic name="inputBitWidth" value="32" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="0.00694153160147458,0.004442905573082777,0.00542809612648147,0.006192842641356624,0.006618294828050123,0.006603562499993257,0.006079175224702046,0.005018467352547563,0.0034449065638808216,0.0014341735004338814,-8.89498572338419E-4,-0.0033627332138082603,-0.005797311285611762,-0.007998295658160745,-0.009783644172042626,-0.011003285120726247,-0.011555421935510976,-0.011398019269542344,-0.010553992198327405,-0.009109275155624125,-0.007204322929741159,-0.005019140044071519,-0.0027540568810415665,-6.083980089812204E-4,0.0012404610374846278,0.0026556133435476385,0.0035540269495699522,0.003913466581767856,0.00377230466955208,0.0032225140769348275,0.0023959414208260354,0.001446970164514328,5.326652362764596E-4,-2.066007958254735E-4,-6.638380285783963E-4,-7.768196094429652E-4,-5.340476658701047E-4,2.62514104027026E-5,8.238895610837434E-4,0.0017486581946731122,0.0026765844956934282,0.003487098913745979,0.004078393178639567,0.00438083982744986,0.0043646125619280045,0.004042076482564693,0.0034650491588244714,0.0027153598060096597,0.0018936995696088965,0.0011044052248033974,4.419334308560773E-4,-2.198853748571485E-5,-2.468668494210699E-4,-2.2794614168577095E-4,4.864160614318245E-6,3.925649504614233E-4,8.56566822210587E-4,0.0013105470106409092,0.0016729586727682298,0.0018782766186860372,0.0018857889745059258,0.0016843460253365488,0.0012928525062685951,7.56475472821023E-4,1.3936353286317209E-4,-4.8498381202610367E-4,-0.0010443810121045153,-0.0014779220044028579,-0.0017442622260908892,-0.0018266948166025957,-0.0017345984228362553,-0.0015011320854918199,-0.0011776820641613787,-8.256332535726899E-4,-5.073585492368197E-4,-2.767953533801635E-4,-1.7243547852371186E-4,-2.116113678975511E-4,-3.9002131744076497E-4,-6.819220738493828E-4,-0.001046019223239551,-0.0014309626704771853,-0.0017834051061336523,-0.002055896030651698,-0.0022127151722109717,-0.002235386631667041,-0.00212450653857447,-0.0018988593120224993,-0.001592730018942093,-0.0012497544795875926,-9.161212222771753E-4,-6.340025728279222E-4,-4.353319446788731E-4,-3.379245812691778E-4,-3.4391279121006614E-4,-4.402790752048672E-4,-6.009333472664914E-4,-7.911330242238177E-4,-9.723698267409983E-4,-0.001108118868193801,-0.001169605167804924,-0.0011403116218206483,-0.0010177282218501317,-8.126308257367965E-4,-5.463585744960325E-4,-2.472163917648406E-4,5.326151816736071E-5,3.236588080786032E-4,5.371302313771076E-4,6.762732858398476E-4,7.365512915308453E-4,7.257403160421124E-4,6.599159361149952E-4,5.595184770490192E-4,4.4835851657187544E-4,3.5356798656509416E-4,3.0020046590606355E-4,3.016124251845741E-4,3.578036877728094E-4,4.6655352894720844E-4,6.249376391672456E-4,8.09643744694843E-4,9.893092489544578E-4,0.0011667674814811555,0.001299313169292976,0.0013897641043404691,0.0014240110405581948,0.0014049635212013609,0.0013390189697002877,0.0012385240475804849,0.001118973010790387,9.968049228555641E-4,8.871151566153326E-4,8.017586589859504E-4,7.479534854997311E-4,7.277751423746349E-4,7.381809738652977E-4,7.717851681733942E-4,8.181696290661348E-4,8.655271963091744E-4,9.021790021476263E-4,9.179025048962746E-4,9.053094830454813E-4,8.604059954823273E-4,7.828479739502213E-4,6.757459764477602E-4,5.452550069508809E-4,3.996345047825579E-4,2.4835564441883347E-4,1.0107320830456308E-4,-3.346298045073322E-5,-1.4841230094082646E-4,-2.3908754151861708E-4,-3.0371511151496537E-4,-3.4334936483498905E-4,-3.6183167642036195E-4,-3.6521146966575225E-4,-3.6143074020422223E-4,-3.590937786685034E-4,-3.667603294346121E-4,-3.921495514277598E-4,-4.4063778119139674E-4,-5.14912732400436E-4,-6.141975134298923E-4,-7.339067709041872E-4,-8.665176616632279E-4,-0.001001720273097524,-0.0011278561006899076,-0.0012334371144421788,-0.00130809901249336,-0.001344930606628321,-0.0013407133554578044,-0.0012973317325593388,-0.0012213045533098353,-0.0011236109470494275,-0.0010181201710717268,-9.200391409651332E-4,-8.4354927594562E-4,-7.996912659978402E-4,-7.945917150000017E-4,-8.283340180089673E-4,-8.945858428943827E-4,-9.813107758859648E-4,-0.00107208268060287,-0.0011483301356481727,-0.0011919580492424074,-0.0011881375908154156,-0.0011277356530553844,-0.0010090479403760733,-8.38590375927257E-4,-6.304185083571683E-4,-4.0444785055313763E-4,-1.836568081101106E-4,9.253774178457668E-6,1.5524828022499458E-4,2.4175987099524617E-4,2.6500500663536144E-4,2.3064997300615252E-4,1.5383076383671635E-4,5.645058414963538E-5,-3.471970902365569E-5,-9.387108763138222E-5,-9.824531544629252E-5,-3.374445743930996E-5,1.0401203059689652E-4,3.082432776944931E-4,5.610392196281046E-4,8.36640113533579E-4,0.0011039575740735541,0.0013313356166386354,0.0014921823309014307,0.001568535651816849,0.0015544366520768933,0.0014572370031299814,0.0012961630417673595,0.0010999602158623626,9.032430599554325E-4,7.412565864967927E-4,6.439479728900315E-4,6.313377834476423E-4,7.096929109839254E-4,8.704050889764356E-4,0.0010913329134503264,0.0013398459419653574,0.0015767722401159806,0.0017621606138371261,0.0018621389621410382,0.0018548888554187693,0.0017338533156117917,0.0015086227022526218,0.0012037818304989926,8.565414847908129E-4,5.116352966694704E-4,2.1364580287916904E-4,-8.253514513628299E-7,-1.0782815677833513E-4,-9.866245104334945E-5,1.6742292393230376E-5,2.0929463820690175E-4,4.3731123462308557E-4,6.544761262929614E-4,8.125814400234609E-4,8.691887206770601E-4,8.010970820737466E-4,6.019243225970459E-4,2.807636322644865E-4,-1.2406504053271455E-4,-5.715091327864377E-4,-0.001003849276949346,-0.001369811050370319,-0.0016242154292971677,-0.0017390327665658752,-0.0017065857370787542,-0.0015416722388411268,-0.0012795551764417403,-9.708260034813308E-4,-6.737215141541751E-4,-4.452935866955523E-4,-3.323464401497307E-4,-3.6378938405269736E-4,-5.456477803203586E-4,-8.597433921520448E-4,-0.001265928273657488,-0.0017077910943735473,-0.0021212041115907954,-0.0024439775446284603,-0.002625691979158311,-0.002635826849854234,-0.0024690173500713612,-0.0021462170070841702,-0.0017120593027541904,-0.001228404584847254,-7.649680691170891E-4,-3.8848678557078914E-4,-1.524511657747846E-4,-8.812526021861288E-5,-1.9959514595421532E-4,-4.6246874820432424E-4,-8.273476247954973E-4,-0.001226718164426176,-0.0015856331100504546,-0.0018330232241552346,-0.001913088073656218,-0.0017947161677516054,-0.0014763758727295226,-9.873982555801857E-4,-3.8393616217254534E-4,2.594805526414807E-4,8.60661129831961E-4,0.00134292120948244,0.0016469102615186944,0.001739984743766607,0.001622302345617116,0.0013266253252058983,9.144282747346136E-4,4.6617856173256886E-4,6.935217790709078E-5,-1.9561085022019176E-4,-2.6783617015077566E-4,-1.1624385929286545E-4,2.550904211323507E-4,8.067919775201523E-4,0.0014695268603228857,0.002154172192559708,0.0027654758798047394,0.0032167396284371015,0.003443680949206284,0.0034148427939363147,0.003137092698585297,0.0026551222581965195,0.0020451537620904217,0.0014036254069544542,8.323369966807399E-4,4.226681183004021E-4,2.4087606728696176E-4,3.1711376935072977E-4,6.399951266359329E-4,0.0011577434769828754,0.0017854744325133444,0.0024180946100370495,0.0029460094792129014,0.003272879570541053,0.003329873519540327,0.0030891566035878503,0.0025664853292876174,0.0018225733364971234,9.515244953826791E-4,6.861907247022276E-5,-7.075147311377331E-4,-0.0012743854126327846,-0.001560419486337564,-0.0015378599531795034,-0.0012282145041799526,-6.985151746065434E-4,-5.22672580313851E-5,5.860813735181133E-4,0.0010908930315750214,0.0013547634109130765,0.0013057710082329662,9.202482401364109E-4,2.276276610249278E-4,-6.939261418451777E-4,-0.0017283413549499247,-0.0027385896670985956,-0.003587666499137697,-0.004160539191487493,-0.004382525797213568,-0.004231582036492468,-0.003742549505946583,-0.003002842779247927,-0.002139895374015729,-0.0013019924310194823,-6.34649653799084E-4,-2.5761571403982357E-4,-2.458628129200586E-4,-6.169201023451345E-4,-0.001325901633780712,-0.002271369980453547,-0.003311116137677649,-0.004282972978415425,-0.005028826507403592,-0.005420924664105858,-0.005383442173331444,-0.004903052560735484,-0.004033473481675513,-0.0028910093497948202,-0.0016336023381956304,-4.385329721366788E-4,5.218853923734076E-4,0.0011149354463698418,0.0012599904351450414,9.508314559172937E-4,2.522664204699066E-4,-7.048504661279154E-4,-0.00174476100158851,-0.0026726719161245514,-0.0033053407814170395,-0.0035002808227615656,-0.0031795406358179268,-0.0023436911974200137,-0.0010738736211853854,4.7886433620265785E-4,0.0021154294660078645,0.0036187242566496267,0.004787058994938294,0.005466231587808179,0.005575094831076192,0.005120019313220455,0.004196097330928216,0.002974278143108524,0.0016763722388929267,5.411835859467459E-4,-2.127117219768144E-4,-4.2225582639876806E-4,-7.50137255929945E-6,0.0010131821681000008,0.002523136823771827,0.004322427479081041,0.006157021796823805,0.007756741472285695,0.008877485809280716,0.009340075158046704,0.00906091815113947,0.008067566669650243,0.006498080088340594,0.004582753410074113,0.0026103819422979018,8.851206256911547E-4,-3.214309269387653E-4,-8.142678074038249E-4,-5.08208413543875E-4,5.541957414329669E-4,0.002205199786489506,0.004173585776594425,0.006123303471739178,0.007704486645810512,0.008607433569503562,0.008613551867194343,0.007633137395800894,0.005725139544675453,0.0030937517627687315,6.270487071321271E-5,-0.0029707748346615094,-0.005595097083141493,-0.007448236106760472,-0.008276787051412366,-0.007980803835215135,-0.006636548240081061,-0.0044930446031293475,-0.001941243656435793,5.403814220775672E-4,0.0024566717032864405,0.003372604567429888,0.0029849261732649976,0.001177308764045355,-0.0019505736410855,-0.006085512406536623,-0.010736516170794519,-0.015300079266471905,-0.019146669264065733,-0.021716327426916506,-0.022610028253282084,-0.021662256644977843,-0.01898378613946548,-0.014963991419854666,-0.010234512627906091,-0.005588625171058915,-0.0018784451464396552,1.1409649234494087E-4,-2.0341741963661637E-4,-0.003124937506393118,-0.008573131850591564,-0.016075194147092273,-0.02478694164235587,-0.03357210887303145,-0.04112715010294271,-0.046134539979822045,-0.04743078468693403,-0.04416671187991793,-0.035936516234332694,-0.022859655139752764,-0.005604352318506481,0.014654476575978823,0.03634052422327449,0.05763186436790323,0.07665074179381524,0.09166538248916777,0.10128000332779885,0.10458937104329608,0.10128000332779885,0.09166538248916777,0.07665074179381524,0.05763186436790323,0.03634052422327449,0.014654476575978823,-0.005604352318506481,-0.022859655139752764,-0.035936516234332694,-0.04416671187991793,-0.04743078468693403,-0.046134539979822045,-0.04112715010294271,-0.03357210887303145,-0.02478694164235587,-0.016075194147092273,-0.008573131850591564,-0.003124937506393118,-2.0341741963661637E-4,1.1409649234494087E-4,-0.0018784451464396552,-0.005588625171058915,-0.010234512627906091,-0.014963991419854666,-0.01898378613946548,-0.021662256644977843,-0.022610028253282084,-0.021716327426916506,-0.019146669264065733,-0.015300079266471905,-0.010736516170794519,-0.006085512406536623,-0.0019505736410855,0.001177308764045355,0.0029849261732649976,0.003372604567429888,0.0024566717032864405,5.403814220775672E-4,-0.001941243656435793,-0.0044930446031293475,-0.006636548240081061,-0.007980803835215135,-0.008276787051412366,-0.007448236106760472,-0.005595097083141493,-0.0029707748346615094,6.270487071321271E-5,0.0030937517627687315,0.005725139544675453,0.007633137395800894,0.008613551867194343,0.008607433569503562,0.007704486645810512,0.006123303471739178,0.004173585776594425,0.002205199786489506,5.541957414329669E-4,-5.08208413543875E-4,-8.142678074038249E-4,-3.214309269387653E-4,8.851206256911547E-4,0.0026103819422979018,0.004582753410074113,0.006498080088340594,0.008067566669650243,0.00906091815113947,0.009340075158046704,0.008877485809280716,0.007756741472285695,0.006157021796823805,0.004322427479081041,0.002523136823771827,0.0010131821681000008,-7.50137255929945E-6,-4.2225582639876806E-4,-2.127117219768144E-4,5.411835859467459E-4,0.0016763722388929267,0.002974278143108524,0.004196097330928216,0.005120019313220455,0.005575094831076192,0.005466231587808179,0.004787058994938294,0.0036187242566496267,0.0021154294660078645,4.7886433620265785E-4,-0.0010738736211853854,-0.0023436911974200137,-0.0031795406358179268,-0.0035002808227615656,-0.0033053407814170395,-0.0026726719161245514,-0.00174476100158851,-7.048504661279154E-4,2.522664204699066E-4,9.508314559172937E-4,0.0012599904351450414,0.0011149354463698418,5.218853923734076E-4,-4.385329721366788E-4,-0.0016336023381956304,-0.0028910093497948202,-0.004033473481675513,-0.004903052560735484,-0.005383442173331444,-0.005420924664105858,-0.005028826507403592,-0.004282972978415425,-0.003311116137677649,-0.002271369980453547,-0.001325901633780712,-6.169201023451345E-4,-2.458628129200586E-4,-2.5761571403982357E-4,-6.34649653799084E-4,-0.0013019924310194823,-0.002139895374015729,-0.003002842779247927,-0.003742549505946583,-0.004231582036492468,-0.004382525797213568,-0.004160539191487493,-0.003587666499137697,-0.0027385896670985956,-0.0017283413549499247,-6.939261418451777E-4,2.276276610249278E-4,9.202482401364109E-4,0.0013057710082329662,0.0013547634109130765,0.0010908930315750214,5.860813735181133E-4,-5.22672580313851E-5,-6.985151746065434E-4,-0.0012282145041799526,-0.0015378599531795034,-0.001560419486337564,-0.0012743854126327846,-7.075147311377331E-4,6.861907247022276E-5,9.515244953826791E-4,0.0018225733364971234,0.0025664853292876174,0.0030891566035878503,0.003329873519540327,0.003272879570541053,0.0029460094792129014,0.0024180946100370495,0.0017854744325133444,0.0011577434769828754,6.399951266359329E-4,3.1711376935072977E-4,2.4087606728696176E-4,4.226681183004021E-4,8.323369966807399E-4,0.0014036254069544542,0.0020451537620904217,0.0026551222581965195,0.003137092698585297,0.0034148427939363147,0.003443680949206284,0.0032167396284371015,0.0027654758798047394,0.002154172192559708,0.0014695268603228857,8.067919775201523E-4,2.550904211323507E-4,-1.1624385929286545E-4,-2.6783617015077566E-4,-1.9561085022019176E-4,6.935217790709078E-5,4.6617856173256886E-4,9.144282747346136E-4,0.0013266253252058983,0.001622302345617116,0.001739984743766607,0.0016469102615186944,0.00134292120948244,8.60661129831961E-4,2.594805526414807E-4,-3.8393616217254534E-4,-9.873982555801857E-4,-0.0014763758727295226,-0.0017947161677516054,-0.001913088073656218,-0.0018330232241552346,-0.0015856331100504546,-0.001226718164426176,-8.273476247954973E-4,-4.6246874820432424E-4,-1.9959514595421532E-4,-8.812526021861288E-5,-1.524511657747846E-4,-3.8848678557078914E-4,-7.649680691170891E-4,-0.001228404584847254,-0.0017120593027541904,-0.0021462170070841702,-0.0024690173500713612,-0.002635826849854234,-0.002625691979158311,-0.0024439775446284603,-0.0021212041115907954,-0.0017077910943735473,-0.001265928273657488,-8.597433921520448E-4,-5.456477803203586E-4,-3.6378938405269736E-4,-3.323464401497307E-4,-4.452935866955523E-4,-6.737215141541751E-4,-9.708260034813308E-4,-0.0012795551764417403,-0.0015416722388411268,-0.0017065857370787542,-0.0017390327665658752,-0.0016242154292971677,-0.001369811050370319,-0.001003849276949346,-5.715091327864377E-4,-1.2406504053271455E-4,2.807636322644865E-4,6.019243225970459E-4,8.010970820737466E-4,8.691887206770601E-4,8.125814400234609E-4,6.544761262929614E-4,4.3731123462308557E-4,2.0929463820690175E-4,1.6742292393230376E-5,-9.866245104334945E-5,-1.0782815677833513E-4,-8.253514513628299E-7,2.1364580287916904E-4,5.116352966694704E-4,8.565414847908129E-4,0.0012037818304989926,0.0015086227022526218,0.0017338533156117917,0.0018548888554187693,0.0018621389621410382,0.0017621606138371261,0.0015767722401159806,0.0013398459419653574,0.0010913329134503264,8.704050889764356E-4,7.096929109839254E-4,6.313377834476423E-4,6.439479728900315E-4,7.412565864967927E-4,9.032430599554325E-4,0.0010999602158623626,0.0012961630417673595,0.0014572370031299814,0.0015544366520768933,0.001568535651816849,0.0014921823309014307,0.0013313356166386354,0.0011039575740735541,8.36640113533579E-4,5.610392196281046E-4,3.082432776944931E-4,1.0401203059689652E-4,-3.374445743930996E-5,-9.824531544629252E-5,-9.387108763138222E-5,-3.471970902365569E-5,5.645058414963538E-5,1.5383076383671635E-4,2.3064997300615252E-4,2.6500500663536144E-4,2.4175987099524617E-4,1.5524828022499458E-4,9.253774178457668E-6,-1.836568081101106E-4,-4.0444785055313763E-4,-6.304185083571683E-4,-8.38590375927257E-4,-0.0010090479403760733,-0.0011277356530553844,-0.0011881375908154156,-0.0011919580492424074,-0.0011483301356481727,-0.00107208268060287,-9.813107758859648E-4,-8.945858428943827E-4,-8.283340180089673E-4,-7.945917150000017E-4,-7.996912659978402E-4,-8.4354927594562E-4,-9.200391409651332E-4,-0.0010181201710717268,-0.0011236109470494275,-0.0012213045533098353,-0.0012973317325593388,-0.0013407133554578044,-0.001344930606628321,-0.00130809901249336,-0.0012334371144421788,-0.0011278561006899076,-0.001001720273097524,-8.665176616632279E-4,-7.339067709041872E-4,-6.141975134298923E-4,-5.14912732400436E-4,-4.4063778119139674E-4,-3.921495514277598E-4,-3.667603294346121E-4,-3.590937786685034E-4,-3.6143074020422223E-4,-3.6521146966575225E-4,-3.6183167642036195E-4,-3.4334936483498905E-4,-3.0371511151496537E-4,-2.3908754151861708E-4,-1.4841230094082646E-4,-3.346298045073322E-5,1.0107320830456308E-4,2.4835564441883347E-4,3.996345047825579E-4,5.452550069508809E-4,6.757459764477602E-4,7.828479739502213E-4,8.604059954823273E-4,9.053094830454813E-4,9.179025048962746E-4,9.021790021476263E-4,8.655271963091744E-4,8.181696290661348E-4,7.717851681733942E-4,7.381809738652977E-4,7.277751423746349E-4,7.479534854997311E-4,8.017586589859504E-4,8.871151566153326E-4,9.968049228555641E-4,0.001118973010790387,0.0012385240475804849,0.0013390189697002877,0.0014049635212013609,0.0014240110405581948,0.0013897641043404691,0.001299313169292976,0.0011667674814811555,9.893092489544578E-4,8.09643744694843E-4,6.249376391672456E-4,4.6655352894720844E-4,3.578036877728094E-4,3.016124251845741E-4,3.0020046590606355E-4,3.5356798656509416E-4,4.4835851657187544E-4,5.595184770490192E-4,6.599159361149952E-4,7.257403160421124E-4,7.365512915308453E-4,6.762732858398476E-4,5.371302313771076E-4,3.236588080786032E-4,5.326151816736071E-5,-2.472163917648406E-4,-5.463585744960325E-4,-8.126308257367965E-4,-0.0010177282218501317,-0.0011403116218206483,-0.001169605167804924,-0.001108118868193801,-9.723698267409983E-4,-7.911330242238177E-4,-6.009333472664914E-4,-4.402790752048672E-4,-3.4391279121006614E-4,-3.379245812691778E-4,-4.353319446788731E-4,-6.340025728279222E-4,-9.161212222771753E-4,-0.0012497544795875926,-0.001592730018942093,-0.0018988593120224993,-0.00212450653857447,-0.002235386631667041,-0.0022127151722109717,-0.002055896030651698,-0.0017834051061336523,-0.0014309626704771853,-0.001046019223239551,-6.819220738493828E-4,-3.9002131744076497E-4,-2.116113678975511E-4,-1.7243547852371186E-4,-2.767953533801635E-4,-5.073585492368197E-4,-8.256332535726899E-4,-0.0011776820641613787,-0.0015011320854918199,-0.0017345984228362553,-0.0018266948166025957,-0.0017442622260908892,-0.0014779220044028579,-0.0010443810121045153,-4.8498381202610367E-4,1.3936353286317209E-4,7.56475472821023E-4,0.0012928525062685951,0.0016843460253365488,0.0018857889745059258,0.0018782766186860372,0.0016729586727682298,0.0013105470106409092,8.56566822210587E-4,3.925649504614233E-4,4.864160614318245E-6,-2.2794614168577095E-4,-2.468668494210699E-4,-2.198853748571485E-5,4.419334308560773E-4,0.0011044052248033974,0.0018936995696088965,0.0027153598060096597,0.0034650491588244714,0.004042076482564693,0.0043646125619280045,0.00438083982744986,0.004078393178639567,0.003487098913745979,0.0026765844956934282,0.0017486581946731122,8.238895610837434E-4,2.62514104027026E-5,-5.340476658701047E-4,-7.768196094429652E-4,-6.638380285783963E-4,-2.066007958254735E-4,5.326652362764596E-4,0.001446970164514328,0.0023959414208260354,0.0032225140769348275,0.00377230466955208,0.003913466581767856,0.0035540269495699522,0.0026556133435476385,0.0012404610374846278,-6.083980089812204E-4,-0.0027540568810415665,-0.005019140044071519,-0.007204322929741159,-0.009109275155624125,-0.010553992198327405,-0.011398019269542344,-0.011555421935510976,-0.011003285120726247,-0.009783644172042626,-0.007998295658160745,-0.005797311285611762,-0.0033627332138082603,-8.89498572338419E-4,0.0014341735004338814,0.0034449065638808216,0.005018467352547563,0.006079175224702046,0.006603562499993257,0.006618294828050123,0.006192842641356624,0.00542809612648147,0.004442905573082777,0.00694153160147458" />
// Retrieval info: 	<generic name="coeffSetRealValueImag" value="0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, -0.0530093, -0.04498, 0.0, 0.0749693, 0.159034, 0.224907, 0.249809, 0.224907, 0.159034, 0.0749693, 0.0, -0.04498, -0.0530093, -0.0321283, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0" />
// Retrieval info: 	<generic name="coeffScaling" value="auto" />
// Retrieval info: 	<generic name="coeffType" value="int" />
// Retrieval info: 	<generic name="coeffBitWidth" value="10" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffComplex" value="false" />
// Retrieval info: 	<generic name="karatsuba" value="false" />
// Retrieval info: 	<generic name="outType" value="int" />
// Retrieval info: 	<generic name="outMSBRound" value="sat" />
// Retrieval info: 	<generic name="outMsbBitRem" value="20" />
// Retrieval info: 	<generic name="outLSBRound" value="trunc" />
// Retrieval info: 	<generic name="outLsbBitRem" value="0" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : BandFIR5503000.vo
// RELATED_FILES: BandFIR5503000.v, dspba_library_package.vhd, dspba_library.vhd, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, altera_avalon_sc_fifo.v, BandFIR5503000_0002_rtl_core.vhd, BandFIR5503000_0002_ast.vhd, BandFIR5503000_0002.vhd
